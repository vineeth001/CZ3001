library verilog;
use verilog.vl_types.all;
entity alu_tb_file_io is
end alu_tb_file_io;
